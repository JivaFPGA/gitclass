module fa(a, b, c);
endmodule
