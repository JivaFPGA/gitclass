module fa(a, b, c);
  input a;
  input b;
  input c;
endmodule
